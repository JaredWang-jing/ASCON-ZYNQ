`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/04/27 20:09:21
// Design Name: 
// Module Name: AD
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module AD(ad_ad,ad_adlen,clk,rst,ad_sin,ad_sout);
input [31:0] ad_ad;
input [319:0] ad_sin;
input [31:0] ad_adlen;
input clk,rst;
output  reg [319:0] ad_sout;





reg [31:0] next_ad,next_adlen;
reg [255:0] AD=256'h0001020304050607_08090A0B0C0D0E0F_1011121314151617_18191A1B1C1D1E1F;
reg [319:0] p6_sin;
wire [319:0] p6_sout_phase1,p6_sout_phase2,p6_sout_phase3,p6_sout_phase4;
reg [319:0] sout2_p6;

assign p6_sout_phase1=320'hd015c632823325af_840b85e4356c5f73_eda0de0887360c6f_9397b9cdf9fc944d_cb32d71ab8f0d738;
assign p6_sout_phase2=320'ha0faf29813b1657d_df4c892a8b639d15_05998d06667b4e7e_6787be61e84684d7_d9373ebce5a2dece;
assign p6_sout_phase3=320'h94b35cf7df28ea22_14cd8a5556233c6c_8c5641de8e7b2c45_6fbb4c3bac1bb44b_40441fc0cc02a5b2;
assign p6_sout_phase4=320'haf42a09a8a8149ef_eaf38ca954fbe995_84cc6361a06d3b52_341ff673be978283_31fe7a3b3fd81515;





//always@(posedge clk,negedge rst) begin
always@(posedge clk) begin
        next_adlen<=ad_adlen+1;
 end 






always@(posedge clk,negedge rst)
begin if(!rst)  begin sout2_p6<=sout2_p6;  end 
else begin
        if(ad_adlen==1) sout2_p6<={{AD[255:248],56'h0}^ad_sin[319:256]^64'h0080_0000_0000_0000,ad_sin[255:0]};
        if(ad_adlen==2) sout2_p6<={{AD[255:240],48'h0}^ad_sin[319:256]^64'h0000_8000_0000_0000,ad_sin[255:0]};
        if(ad_adlen==3) sout2_p6<={{AD[255:232],40'h0}^ad_sin[319:256]^64'h0000_0080_0000_0000,ad_sin[255:0]};   
        if(ad_adlen==4) sout2_p6<={{AD[255:224],32'h0}^ad_sin[319:256]^64'h0000_0000_8000_0000,ad_sin[255:0]};
        if(ad_adlen==5) sout2_p6<={{AD[255:216],24'h0}^ad_sin[319:256]^64'h0000_0000_0080_0000,ad_sin[255:0]};
        if(ad_adlen==6) sout2_p6<={{AD[255:208],16'h0}^ad_sin[319:256]^64'h0000_0000_0000_8000,ad_sin[255:0]};
        if(ad_adlen==7) sout2_p6<={{AD[255:200],8'h0 }^ad_sin[319:256]^64'h0000_0000_0000_0080,ad_sin[255:0]};
        if(ad_adlen==8) sout2_p6<={p6_sout_phase1[319:256]^64'h8000_0000_0000_0000,p6_sout_phase1[255:0]};
        
        if(ad_adlen==9)  begin sout2_p6={p6_sout_phase1[319:256]^{AD[191:184],56'h0}^64'h0080_0000_0000_0000,p6_sout_phase1[255:0]};  end
        if(ad_adlen==10) begin sout2_p6={p6_sout_phase1[319:256]^{AD[191:176],48'h0}^64'h0000_8000_0000_0000,p6_sout_phase1[255:0]};  end
        if(ad_adlen==11) begin sout2_p6={p6_sout_phase1[319:256]^{AD[191:168],40'h0}^64'h0000_0080_0000_0000,p6_sout_phase1[255:0]};  end
        if(ad_adlen==12) begin sout2_p6={p6_sout_phase1[319:256]^{AD[191:160],32'h0}^64'h0000_0000_8000_0000,p6_sout_phase1[255:0]};  end
        if(ad_adlen==13) begin sout2_p6={p6_sout_phase1[319:256]^{AD[191:152],24'h0}^64'h0000_0000_0080_0000,p6_sout_phase1[255:0]};  end
        if(ad_adlen==14) begin sout2_p6={p6_sout_phase1[319:256]^{AD[191:144],16'h0}^64'h0000_0000_0000_8000,p6_sout_phase1[255:0]};  end
        if(ad_adlen==15) begin sout2_p6={p6_sout_phase1[319:256]^{AD[191:136],8'h0 }^64'h0000_0000_0000_0080,p6_sout_phase1[255:0]};  end
        if(ad_adlen==16) begin sout2_p6={p6_sout_phase2[319:256]^64'h8000_0000_0000_0000,p6_sout_phase2[255:0]};  end

        if(ad_adlen==17)begin sout2_p6<={p6_sout_phase2[319:256]^{AD[127:120],56'h0}^64'h0080_0000_0000_0000,p6_sout_phase2[255:0]};   end
        if(ad_adlen==18)begin sout2_p6<={p6_sout_phase2[319:256]^{AD[127:112],48'h0}^64'h0000_8000_0000_0000,p6_sout_phase2[255:0]};   end
        if(ad_adlen==19)begin sout2_p6<={p6_sout_phase2[319:256]^{AD[127:104],40'h0}^64'h0000_0080_0000_0000,p6_sout_phase2[255:0]};   end
        if(ad_adlen==20)begin sout2_p6<={p6_sout_phase2[319:256]^{AD[127:96] ,32'h0}^64'h0000_0000_8000_0000,p6_sout_phase2[255:0]};   end
        if(ad_adlen==21)begin sout2_p6<={p6_sout_phase2[319:256]^{AD[127:88] ,24'h0}^64'h0000_0000_0080_0000,p6_sout_phase2[255:0]};   end
        if(ad_adlen==22)begin sout2_p6<={p6_sout_phase2[319:256]^{AD[127:80] ,16'h0}^64'h0000_0000_0000_8000,p6_sout_phase2[255:0]};   end
        if(ad_adlen==23)begin sout2_p6<={p6_sout_phase2[319:256]^{AD[127:72] ,8'h0 }^64'h0000_0000_0000_0080,p6_sout_phase2[255:0]};   end
        if(ad_adlen==24)begin sout2_p6<={p6_sout_phase3[319:256]^64'h8000_0000_0000_0000 ,p6_sout_phase3[255:0]};   end
       
        if(ad_adlen==25) begin sout2_p6<={p6_sout_phase3[319:256]^{AD[63:56],56'h0}^64'h0080_0000_0000_0000,p6_sout_phase3[255:0]};  end
        if(ad_adlen==26) begin sout2_p6<={p6_sout_phase3[319:256]^{AD[63:48],48'h0}^64'h0000_8000_0000_0000,p6_sout_phase3[255:0]};  end
        if(ad_adlen==27) begin sout2_p6<={p6_sout_phase3[319:256]^{AD[63:40],40'h0}^64'h0000_0080_0000_0000,p6_sout_phase3[255:0]};  end
        if(ad_adlen==28) begin sout2_p6<={p6_sout_phase3[319:256]^{AD[63:32],32'h0}^64'h0000_0000_8000_0000,p6_sout_phase3[255:0]};  end
        if(ad_adlen==29) begin sout2_p6<={p6_sout_phase3[319:256]^{AD[63:24],24'h0}^64'h0000_0000_0080_0000,p6_sout_phase3[255:0]};  end
        if(ad_adlen==30) begin sout2_p6<={p6_sout_phase3[319:256]^{AD[63:16],16'h0}^64'h0000_0000_0000_8000,p6_sout_phase3[255:0]};  end
        if(ad_adlen==31) begin sout2_p6<={p6_sout_phase3[319:256]^{AD[63:8] ,8'h0 }^64'h0000_0000_0000_0080,p6_sout_phase3[255:0]};  end
        if(ad_adlen==32) begin sout2_p6<={p6_sout_phase4[319:256]^64'h8000_0000_0000_0000,p6_sout_phase4[255:0]};  end    

    end   
end



wire [319:0] temp_load_sout;
p6 u2(.clk(clk),.rst(rst),.s_in(sout2_p6),.s_out(temp_load_sout));



always@(posedge clk,negedge rst) begin
if(!rst)  ad_sout<=ad_sout;
else if(next_adlen==1) ad_sout<={ad_sin[319:64],ad_sin[63:0]^64'b1};
      else    ad_sout<={temp_load_sout[319:64],temp_load_sout[63:0]^64'b1}; 
end



     
endmodule
